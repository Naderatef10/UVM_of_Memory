package pack1;

import uvm_pkg::*;


`include "uvm_macros.svh"

`include "interface.sv"
`include "low_sequence_item.sv"
`include "low_sequencer.sv"
`include "low_driver.sv"
`include "low_monitor.sv"

`include "low_agent.sv"
`include "low_scoreboard.sv"
`include "low_subscriber.sv"

`include "low_env.sv"
`include "low_test.sv"

endpackage

